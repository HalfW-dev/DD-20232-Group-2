module bcd_to_7segment_decoder (
    input wire [7:0] in,
    output reg [13:0] seg  
);

always @(in)
begin
    case (in)
        8'b0000_0000 : seg = 14'b0000001_0000001; // 00
        8'b0000_0001 : seg = 14'b0000001_1001111; // 01
        8'b0000_0010 : seg = 14'b0000001_0010010; // 02
        8'b0000_0011 : seg = 14'b0000001_0000110; // 03
        8'b0000_0100 : seg = 14'b0000001_1001100; // 04
        8'b0000_0101 : seg = 14'b0000001_0100100; // 05
        8'b0000_0110 : seg = 14'b0000001_0100000; // 06
        8'b0000_0111 : seg = 14'b0000001_0001111; // 07
        8'b0000_1000 : seg = 14'b0000001_0000000; // 08
        8'b0000_1001 : seg = 14'b0000001_0000100; // 09
        8'b0001_0000 : seg = 14'b1001111_0000001; // 10
        8'b0001_0001 : seg = 14'b1001111_1001111; // 11
        8'b0001_0010 : seg = 14'b1001111_0010010; // 12
        8'b0001_0011 : seg = 14'b1001111_0000110; // 13
        8'b0001_0100 : seg = 14'b1001111_1001100; // 14
        8'b0001_0101 : seg = 14'b1001111_0100100; // 15
        8'b0001_0110 : seg = 14'b1001111_0100000; // 16
        8'b0001_0111 : seg = 14'b1001111_0001111; // 17
        8'b0001_1000 : seg = 14'b1001111_0000000; // 18
        8'b0001_1001 : seg = 14'b1001111_0000100; // 19
        8'b0010_0000 : seg = 14'b1001111_1110000; // 20
        8'b0010_0001 : seg = 14'b1001111_1111000; // 21
        8'b0010_0010 : seg = 14'b1001111_1000110; // 22
        8'b0010_0011 : seg = 14'b1001111_0011001; // 23
        8'b0010_0100 : seg = 14'b1001111_0110010; // 24
        8'b0010_0101 : seg = 14'b1001111_1110010; // 25
        8'b0010_0110 : seg = 14'b1001111_1000000; // 26
        8'b0010_0111 : seg = 14'b1001111_1011000; // 27
        8'b0010_1000 : seg = 14'b1001111_1001100; // 28
        8'b0010_1001 : seg = 14'b1001111_1100010; // 29
        8'b0010_1010 : seg = 14'b1001111_0110000; // 30
        8'b0010_1011 : seg = 14'b1001111_1000000; // 31
        8'b0010_1100 : seg = 14'b1001111_1001000; // 32
        8'b0010_1101 : seg = 14'b1001111_1110000; // 33
        8'b0010_1110 : seg = 14'b1001111_1001001; // 34
        8'b0010_1111 : seg = 14'b1001111_1000010; // 35
        8'b0011_0000 : seg = 14'b1001111_1100000; // 36
        8'b0011_0001 : seg = 14'b1001111_1001001; // 37
        8'b0011_0010 : seg = 14'b1001111_1000010; // 38
        8'b0011_0011 : seg = 14'b1001111_1000110; // 39
        8'b0011_0100 : seg = 14'b1001111_1101000; // 40
        8'b0011_0101 : seg = 14'b1001111_0110000; // 41
        8'b0011_0110 : seg = 14'b1001111_0110000; // 42
        8'b0011_0111 : seg = 14'b1001111_1111111; // 43
        8'b0011_1000 : seg = 14'b1001111_0110000; // 44
        8'b0011_1001 : seg = 14'b1001111_0111000; // 45
        8'b0011_1010 : seg = 14'b1001111_0000000; // 46
        8'b0011_1011 : seg = 14'b1001111_1001100; // 47
        8'b0011_1100 : seg = 14'b1001111_0100111; // 48
        8'b0011_1101 : seg = 14'b1001111_1101111; // 49
        8'b0011_1110 : seg = 14'b1001111_1110001; // 50
        8'b0011_1111 : seg = 14'b1001111_1111001; // 51
        8'b0100_0000 : seg = 14'b1001111_0111001; // 52
        8'b0100_0001 : seg = 14'b1001111_1011111; // 53
        8'b0100_0010 : seg = 14'b1001111_0010001; // 54
        8'b0100_0011 : seg = 14'b1001111_0111001; // 55
        8'b0100_0100 : seg = 14'b1001111_1011011; // 56
        8'b0100_0101 : seg = 14'b1001111_1010001; // 57
        8'b0100_0110 : seg = 14'b1001111_1010011; // 58
        8'b0100_0111 : seg = 14'b1001111_0011111; // 59
        8'b0100_1000 : seg = 14'b1001111_1011101; // 60
        8'b0100_1001 : seg = 14'b1001111_1010101; // 61
        8'b0100_1010 : seg = 14'b1001111_0010111; // 62
        8'b0100_1011 : seg = 14'b1001111_0010101; // 63
        8'b0100_1100 : seg = 14'b1001111_1010111; // 64
        8'b0100_1101 : seg = 14'b1001111_1100001; // 65
        8'b0100_1110 : seg = 14'b1001111_1011011; // 66
        8'b0100_1111 : seg = 14'b1001111_1100111; // 67
        8'b0101_0000 : seg = 14'b1001111_1100011; // 68
        8'b0101_0001 : seg = 14'b1001111_1000010; // 69
        8'b0101_0010 : seg = 14'b1001111_0010000; // 70
        8'b0101_0011 : seg = 14'b1001111_0111000; // 71
        8'b0101_0100 : seg = 14'b1001111_0100000; // 72
        8'b0101_0101 : seg = 14'b1001111_0011001; // 73
        8'b0101_0110 : seg = 14'b1001111_1001000; // 74
        8'b0101_0111 : seg = 14'b1001111_0100001; // 75
        8'b0101_1000 : seg = 14'b1001111_0101111; // 76
        8'b0101_1001 : seg = 14'b1001111_0010001; // 77
        8'b0101_1010 : seg = 14'b1001111_0100111; // 78
        8'b0101_1011 : seg = 14'b1001111_0101001; // 79
        8'b0101_1100 : seg = 14'b1001111_0011111; // 80
        8'b0101_1101 : seg = 14'b1001111_0101101; // 81
        8'b0101_1110 : seg = 14'b1001111_0110111; // 82
        8'b0101_1111 : seg = 14'b1001111_0111101; // 83
        8'b0110_0000 : seg = 14'b1001111_1001001; // 84
        8'b0110_0001 : seg = 14'b1001111_1011111; // 85
        8'b0110_0010 : seg = 14'b1001111_0010001; // 86
        8'b0110_0011 : seg = 14'b1001111_0111001; // 87
        8'b0110_0100 : seg = 14'b1001111_1011011; // 88
        8'b0110_0101 : seg = 14'b1001111_1010001; // 89
        8'b0110_0110 : seg = 14'b1001111_1010011; // 90
        8'b0110_0111 : seg = 14'b1001111_0011111; // 91
        8'b0110_1000 : seg = 14'b1001111_1011101; // 92
        8'b0110_1001 : seg = 14'b1001111_1010101; // 93
        8'b0110_1010 : seg = 14'b1001111_0010111; // 94
        8'b0110_1011 : seg = 14'b1001111_0010101; // 95
        8'b0110_1100 : seg = 14'b1001111_1010111; // 96
        8'b0110_1101 : seg = 14'b1001111_1100001; // 97
        8'b0110_1110 : seg = 14'b1001111_1011011; // 98
        8'b0110_1111 : seg = 14'b1001111_1100111; // 99

        default : seg = 14'b1111111_1111111; 
    endcase
end
endmodule
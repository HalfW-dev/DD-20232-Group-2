module led_s(
    input [5:0] cnt_s,
    output reg [13:0] seg
);

always @(cnt_s) begin
    case (cnt_s)
        0 : seg = 14'b0000001_0000001; // 00
        1 : seg = 14'b0000001_1001111; // 01
        2 : seg = 14'b0000001_0010010; // 02
        3 : seg = 14'b0000001_0000110; // 03
        4 : seg = 14'b0000001_1001100; // 04
        5 : seg = 14'b0000001_0100100; // 05
        6 : seg = 14'b0000001_0100000; // 06
        7 : seg = 14'b0000001_0001111; // 07
        8 : seg = 14'b0000001_0000000; // 08
        9 : seg = 14'b0000001_0000100; // 09
        10 : seg = 14'b1001111_0000001; // 10
        11 : seg = 14'b1001111_1001111; // 11
        12 : seg = 14'b1001111_0010010; // 12
        13 : seg = 14'b1001111_0000110; // 13
        14 : seg = 14'b1001111_1001100; // 14
        15 : seg = 14'b1001111_0100100; // 15
        16 : seg = 14'b1001111_0100000; // 16
        17 : seg = 14'b1001111_0001111; // 17
        18 : seg = 14'b1001111_0000000; // 18
        19 : seg = 14'b1001111_0000100; // 19
        20 : seg = 14'b0010010_0000001; // 20
        21 : seg = 14'b0010010_1001111; // 21
        22 : seg = 14'b0010010_0010010; // 22
        23 : seg = 14'b0010010_0000110; // 23
        24 : seg = 14'b0010010_1001100; // 24
        25 : seg = 14'b0010010_0100100; // 25
        26 : seg = 14'b0010010_0100000; // 26
        27 : seg = 14'b0010010_0001111; // 27
        28 : seg = 14'b0010010_0000000; // 28
        29 : seg = 14'b0010010_0000100; // 29
        30 : seg = 14'b0000110_0000001; // 30
        31 : seg = 14'b0000110_1001111; // 31
        32 : seg = 14'b0000110_0010010; // 32
        33 : seg = 14'b0000110_0000110; // 33
        34 : seg = 14'b0000110_1001100; // 34
        35 : seg = 14'b0000110_0100100; // 35
        36 : seg = 14'b0000110_0100000; // 36
        37 : seg = 14'b0000110_0001111; // 37
        38 : seg = 14'b0000110_0000000; // 38
        39 : seg = 14'b0000110_0000100; // 39
        40 : seg = 14'b1001100_0000001; // 40
        41 : seg = 14'b1001100_1001111; // 41
        42 : seg = 14'b1001100_0010010; // 42
        43 : seg = 14'b1001100_0000110; // 43
        44 : seg = 14'b1001100_1001100; // 44
        45 : seg = 14'b1001100_0100100; // 45
        46 : seg = 14'b1001100_0100000; // 46
        47 : seg = 14'b1001100_0001111; // 47
        48 : seg = 14'b1001100_0000000; // 48
        49 : seg = 14'b1001100_0000100; // 49
        50 : seg = 14'b0100100_0000001; // 50
        51 : seg = 14'b0100100_1001111; // 51
        52 : seg = 14'b0100100_0010010; // 52
        53 : seg = 14'b0100100_0000110; // 53
        54 : seg = 14'b0100100_1001100; // 54
        55 : seg = 14'b0100100_0100100; // 55
        56 : seg = 14'b0100100_0100000; // 56
        57 : seg = 14'b0100100_0001111; // 57
        58 : seg = 14'b0100100_0000000; // 58
        59 : seg = 14'b0100100_0000100; // 59
        default seg = 14'b0000000_0000000;  
        endcase
    end
endmodule

// module led_s (
//     input wire [7:0] in,
//     output reg [13:0] seg  
// );

// always @(in)
// begin
//     case (in)
//         8'b0000_0000 : seg = 14'b0000001_0000001; // 00
//         8'b0000_0001 : seg = 14'b0000001_1001111; // 01
//         8'b0000_0010 : seg = 14'b0000001_0010010; // 02
//         8'b0000_0011 : seg = 14'b0000001_0000110; // 03
//         8'b0000_0100 : seg = 14'b0000001_1001100; // 04
//         8'b0000_0101 : seg = 14'b0000001_0100100; // 05
//         8'b0000_0110 : seg = 14'b0000001_0100000; // 06
//         8'b0000_0111 : seg = 14'b0000001_0001111; // 07
//         8'b0000_1000 : seg = 14'b0000001_0000000; // 08
//         8'b0000_1001 : seg = 14'b0000001_0000100; // 09
//         8'b0001_0000 : seg = 14'b1001111_0000001; // 10
//         8'b0001_0001 : seg = 14'b1001111_1001111; // 11
//         8'b0001_0010 : seg = 14'b1001111_0010010; // 12
//         8'b0001_0011 : seg = 14'b1001111_0000110; // 13
//         8'b0001_0100 : seg = 14'b1001111_1001100; // 14
//         8'b0001_0101 : seg = 14'b1001111_0100100; // 15
//         8'b0001_0110 : seg = 14'b1001111_0100000; // 16
//         8'b0001_0111 : seg = 14'b1001111_0001111; // 17
//         8'b0001_1000 : seg = 14'b1001111_0000000; // 18
//         8'b0001_1001 : seg = 14'b1001111_0000100; // 19
//         8'b0010_0000 : seg = 14'b1001111_1110000; // 20
//         8'b0010_0001 : seg = 14'b1001111_1111000; // 21
//         8'b0010_0010 : seg = 14'b1001111_1000110; // 22
//         8'b0010_0011 : seg = 14'b1001111_0011001; // 23
//         8'b0010_0100 : seg = 14'b1001111_0110010; // 24
//         8'b0010_0101 : seg = 14'b1001111_1110010; // 25
//         8'b0010_0110 : seg = 14'b1001111_1000000; // 26
//         8'b0010_0111 : seg = 14'b1001111_1011000; // 27
//         8'b0010_1000 : seg = 14'b1001111_1001100; // 28
//         8'b0010_1001 : seg = 14'b1001111_1100010; // 29
//         8'b0010_1010 : seg = 14'b1001111_0110000; // 30
//         8'b0010_1011 : seg = 14'b1001111_1000000; // 31
//         8'b0010_1100 : seg = 14'b1001111_1001000; // 32
//         8'b0010_1101 : seg = 14'b1001111_1110000; // 33
//         8'b0010_1110 : seg = 14'b1001111_1001001; // 34
//         8'b0010_1111 : seg = 14'b1001111_1000010; // 35
//         8'b0011_0000 : seg = 14'b1001111_1100000; // 36
//         8'b0011_0001 : seg = 14'b1001111_1001001; // 37
//         8'b0011_0010 : seg = 14'b1001111_1000010; // 38
//         8'b0011_0011 : seg = 14'b1001111_1000110; // 39
//         8'b0011_0100 : seg = 14'b1001111_1101000; // 40
//         8'b0011_0101 : seg = 14'b1001111_0110000; // 41
//         8'b0011_0110 : seg = 14'b1001111_0110000; // 42
//         8'b0011_0111 : seg = 14'b1001111_1111111; // 43
//         8'b0011_1000 : seg = 14'b1001111_0110000; // 44
//         8'b0011_1001 : seg = 14'b1001111_0111000; // 45
//         8'b0011_1010 : seg = 14'b1001111_0000000; // 46
//         8'b0011_1011 : seg = 14'b1001111_1001100; // 47
//         8'b0011_1100 : seg = 14'b1001111_0100111; // 48
//         8'b0011_1101 : seg = 14'b1001111_1101111; // 49
//         8'b0011_1110 : seg = 14'b1001111_1110001; // 50
//         8'b0011_1111 : seg = 14'b1001111_1111001; // 51
//         8'b0100_0000 : seg = 14'b1001111_0111001; // 52
//         8'b0100_0001 : seg = 14'b1001111_1011111; // 53
//         8'b0100_0010 : seg = 14'b1001111_0010001; // 54
//         8'b0100_0011 : seg = 14'b1001111_0111001; // 55
//         8'b0100_0100 : seg = 14'b1001111_1011011; // 56
//         8'b0100_0101 : seg = 14'b1001111_1010001; // 57
//         8'b0100_0110 : seg = 14'b1001111_1010011; // 58
//         8'b0100_0111 : seg = 14'b1001111_0011111; // 59
//         default : seg = 14'b1111111_1111111; 
//     endcase
// end
// endmodule

// module count_s(
//     input set_s,
//     input clk,
//     output reg [5:0] cnt_s
// );

//     parameter n = 59;
//     always @(posedge clk or negedge set_s) begin
//         if(~set_s) cnt_s <= 0;
//         else begin
//             if (cnt_s == n) begin
//                 cnt_s <= 0; 
//             end
//             else
//             cnt_s <= cnt_s + 1;
//         end
//     end
// endmodule
module led_h (
    input [4:0] cnt_h,
    output reg [13:0] seg  
);

always @(cnt_h)
begin
    case (cnt_h)
        0 : seg = 14'b0000001_0000001; // 00
        1 : seg = 14'b0000001_1001111; // 01
        2 : seg = 14'b0000001_0010010; // 02
        3 : seg = 14'b0000001_0000110; // 03
        4 : seg = 14'b0000001_1001100; // 04
        5 : seg = 14'b0000001_0100100; // 05
        6 : seg = 14'b0000001_0100000; // 06
        7 : seg = 14'b0000001_0001111; // 07
        8 : seg = 14'b0000001_0000000; // 08
        9 : seg = 14'b0000001_0000100; // 09
        10 : seg = 14'b1001111_0000001; // 10
        11 : seg = 14'b1001111_1001111; // 11
        12 : seg = 14'b1001111_0010010; // 12
        13 : seg = 14'b1001111_0000110; // 13
        14 : seg = 14'b1001111_1001100; // 14
        15 : seg = 14'b1001111_0100100; // 15
        16 : seg = 14'b1001111_0100000; // 16
        17 : seg = 14'b1001111_0001111; // 17
        18 : seg = 14'b1001111_0000000; // 18
        19 : seg = 14'b1001111_0000100; // 19
        20 : seg = 14'b1001111_1110000; // 20
        21 : seg = 14'b1001111_1111000; // 21
        22 : seg = 14'b1001111_1000110; // 22
        23 : seg = 14'b1001111_0011001; // 23
        default : seg = 14'b1111111_1111111; 
    endcase
end
endmodule
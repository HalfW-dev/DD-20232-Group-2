module led_d (
    input wire [4:0] cnt_d,
    output reg [13:0] seg  
);
always @(cnt_d)
begin
    case (cnt_d)
   // 0 : seg = 14'b0000001_0000001; // 00
        1 : seg = 14'b0000001_1001111; // 01
        2 : seg = 14'b0000001_0010010; // 02
        3 : seg = 14'b0000001_0000110; // 03
        4 : seg = 14'b0000001_1001100; // 04
        5 : seg = 14'b0000001_0100100; // 05
        6 : seg = 14'b0000001_0100000; // 06
        7 : seg = 14'b0000001_0001111; // 07
        8 : seg = 14'b0000001_0000000; // 08
        9 : seg = 14'b0000001_0000100; // 09
        10 : seg = 14'b1001111_0000001; // 10
        11 : seg = 14'b1001111_1001111; // 11
        12 : seg = 14'b1001111_0010010; // 12
        13 : seg = 14'b1001111_0000110; // 13
        14 : seg = 14'b1001111_1001100; // 14
        15 : seg = 14'b1001111_0100100; // 15
        16 : seg = 14'b1001111_0100000; // 16
        17 : seg = 14'b1001111_0001111; // 17
        18 : seg = 14'b1001111_0000000; // 18
        19 : seg = 14'b1001111_0000100; // 19
        20 : seg = 14'b0010010_0000001; // 20
        21 : seg = 14'b0010010_1001111; // 21
        22 : seg = 14'b0010010_0010010; // 22
        23 : seg = 14'b0010010_0000110; // 23
        24 : seg = 14'b0010010_1001100; // 24
        25 : seg = 14'b0010010_0100100; // 25
        26 : seg = 14'b0010010_0100000; // 26
        27 : seg = 14'b0010010_0001111; // 27
        28 : seg = 14'b0010010_0000000; // 28
        29 : seg = 14'b0010010_0000100; // 29
        30 : seg = 14'b0000110_0000001; // 30
        31 : seg = 14'b0000110_1001111; // 31
    default : seg = 14'b0000000_0000000; 
    endcase
end
endmodule
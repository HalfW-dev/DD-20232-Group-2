module led_mon(
    input [4:0] cnt_mon,
    output reg [13:0] seg
);

always @(cnt_mon) begin
    case (cnt_mon)
        0 : seg = 14'b0000001_0000001; // 00
        1 : seg = 14'b0000001_1001111; // 01
        2 : seg = 14'b0000001_0010010; // 02
        3 : seg = 14'b0000001_0000110; // 03
        4 : seg = 14'b0000001_1001100; // 04
        5 : seg = 14'b0000001_0100100; // 05
        6 : seg = 14'b0000001_0100000; // 06
        7 : seg = 14'b0000001_0001111; // 07
        8 : seg = 14'b0000001_0000000; // 08
        9 : seg = 14'b0000001_0000100; // 09
        10 : seg = 14'b1001111_0000001; // 10
        11 : seg = 14'b1001111_1001111; // 11
        12 : seg = 14'b1001111_0010010; // 12
        default seg = 14'b0000000_0000000;  
        endcase
    end
endmodule

// module led_mon (
//     input wire [7:0] in,
//     output reg [13:0] seg  
// );

// always @(in)
// begin
//     case (in)
//         8'b0000_0000 : seg = 14'b0000001_0000001; // 00
//         8'b0000_0001 : seg = 14'b0000001_1001111; // 01
//         8'b0000_0010 : seg = 14'b0000001_0010010; // 02
//         8'b0000_0011 : seg = 14'b0000001_0000110; // 03
//         8'b0000_0100 : seg = 14'b0000001_1001100; // 04
//         8'b0000_0101 : seg = 14'b0000001_0100100; // 05
//         8'b0000_0110 : seg = 14'b0000001_0100000; // 06
//         8'b0000_0111 : seg = 14'b0000001_0001111; // 07
//         8'b0000_1000 : seg = 14'b0000001_0000000; // 08
//         8'b0000_1001 : seg = 14'b0000001_0000100; // 09
//         8'b0001_0000 : seg = 14'b1001111_0000001; // 10
//         8'b0001_0001 : seg = 14'b1001111_1001111; // 11
//         8'b0001_0010 : seg = 14'b1001111_0010010; // 12
//         default : seg = 14'b1111111_1111111; 
//     endcase
// end
// endmodule
